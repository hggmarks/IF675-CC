`timescale 1ms / 1ms
`include "mux_8to1.v"

module mux_8to1_tb;
    wire F;
    reg [7:0] A;
    reg [2:0] Sel;

    mux_8to1_A uut(F, A, Sel);
    mux_8to1_A dut(F, A, Sel);

    initial begin

        $dumpfile("mux_8to1_tb.vcd");
        $dumpvars(0, mux_8to1_tb);

        Sel = 3'b000;    #50;
        A = 8'b00000001; #50;
        A = 8'b00000010; #50;
        A = 8'b00000100; #50;
        A = 8'b00001000; #50;
        A = 8'b00010000; #50;
        A = 8'b00100000; #50;
        A = 8'b01000000; #50;
        A = 8'b10000000; #50;
        A = 8'b00000000;

        Sel = 3'b001;    #50;
        A = 8'b00000001; #50;
        A = 8'b00000010; #50;
        A = 8'b00000100; #50;
        A = 8'b00001000; #50;
        A = 8'b00010000; #50;
        A = 8'b00100000; #50;
        A = 8'b01000000; #50;
        A = 8'b10000000; #50;
        A = 8'b00000000;

        Sel = 3'b010;    #50;
        A = 8'b00000001; #50;
        A = 8'b00000010; #50;
        A = 8'b00000100; #50;
        A = 8'b00001000; #50;
        A = 8'b00010000; #50;
        A = 8'b00100000; #50;
        A = 8'b01000000; #50;
        A = 8'b10000000; #50;
        A = 8'b00000000;

        Sel = 3'b011;    #50;
        A = 8'b00000001; #50;
        A = 8'b00000010; #50;
        A = 8'b00000100; #50;
        A = 8'b00001000; #50;
        A = 8'b00010000; #50;
        A = 8'b00100000; #50;
        A = 8'b01000000; #50;
        A = 8'b10000000; #50;
        A = 8'b00000000;

        Sel = 3'b100;    #50;
        A = 8'b00000001; #50;
        A = 8'b00000010; #50;
        A = 8'b00000100; #50;
        A = 8'b00001000; #50;
        A = 8'b00010000; #50;
        A = 8'b00100000; #50;
        A = 8'b01000000; #50;
        A = 8'b10000000; #50;
        A = 8'b00000000;


        Sel = 3'b101;    #50;
        A = 8'b00000001; #50;
        A = 8'b00000010; #50;
        A = 8'b00000100; #50;
        A = 8'b00001000; #50;
        A = 8'b00010000; #50;
        A = 8'b00100000; #50;
        A = 8'b01000000; #50;
        A = 8'b10000000; #50;
        A = 8'b00000000;

        Sel = 3'b110; #50;
        A = 8'b00000001; #50;
        A = 8'b00000010; #50;
        A = 8'b00000100; #50;
        A = 8'b00001000; #50;
        A = 8'b00010000; #50;
        A = 8'b00100000; #50;
        A = 8'b01000000; #50;
        A = 8'b10000000; #50;
        A = 8'b00000000;


        Sel = 3'b111;    #50;
        A = 8'b00000001; #50;
        A = 8'b00000010; #50;
        A = 8'b00000100; #50;
        A = 8'b00001000; #50;
        A = 8'b00010000; #50;
        A = 8'b00100000; #50;
        A = 8'b01000000; #50;
        A = 8'b10000000; #50;
        A = 8'b00000000;
    end
endmodule

